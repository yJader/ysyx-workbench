module example();
    initial begin $display("Hello World"); $finish; end
endmodule
